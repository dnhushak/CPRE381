-------------------------------------------------------------------------
-- Joseph Zambreno
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- inv.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 1-input NOT 
-- gate.
--
--
-- NOTES:
-- 8/27/08 by JAZ::Design created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity onescomplementer is
  generic(N : integer);
  port(i_A  : in std_logic_vector(N-1 downto 0);
       o_F  : out std_logic_vector(N-1 downto 0));

end onescomplementer;

architecture structure of onescomplementer is

  component inv
    port(i_A             : in std_logic;
         o_F             : out std_logic);
  end component;
  
  
begin
  
    gen_inv: for I in 0 to N-1 generate
      invX : inv 
      port map(i_A => i_A(I),
               o_F => o_F(I));
    end generate gen_inv;
  
end structure;
