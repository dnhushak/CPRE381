-------------------------------------------------------------------------
-- Joseph Zambreno
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- tb_and2.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a simple VHDL testbench for the
-- 2-input AND gate.
--
--
-- NOTES:
-- 8/31/08 by JAZ::Design created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

-- This is an empty entity so we don't need to declare ports
entity onecomptest is

end onecomptest;

architecture behavior of onecomptest is


-- Declare the component we are going to instantiate

component onescomplementer
generic(N : integer := 32);
  port(i_A  : in std_logic_vector(N-1 downto 0);
       o_F  : out std_logic_vector(N-1 downto 0));

end component;

component onescomplementerdataflow
generic(N : integer := 32);
  port(i_A  : in std_logic_vector(N-1 downto 0);
       o_F  : out std_logic_vector(N-1 downto 0));

end component;

-- Signals to connect to the and2 module
signal s_AVector, s_StructVector, S_DataVector: std_logic_vector(31 downto 0);

begin

DUT: onescomplementer
  port map( i_A  => s_AVector,
            o_F  => s_StructVector);
            
DUT2: onescomplementerdataflow
  port map( i_A  => s_AVector,
            o_F  => s_DataVector);

  -- Remember, a process executes sequentially
  -- and then if not told to 'wait' loops back
  -- around
  process
  begin
    s_AVector <= "00000000000000000000000000000000";
    wait for 10 ns;
    
    for I in 0 to 31 loop
      s_AVector(I) <= '1';
      wait for 10 ns;
    end loop;


end process;
end behavior;
